arch aarch64

objects {
cspace_crasher = cnode (8 bits)
cspace_goodbye = cnode (8 bits)
cspace_hello = cnode (8 bits)
cspace_monitor = cnode (8 bits)
frame_crasher_elf_0000 = frame (4k, fill: [{0 768 CDL_FrameFill_FileData "crasher.elf" 65536}])
frame_crasher_elf_0001 = frame (4k, fill: [{0 8 CDL_FrameFill_FileData "crasher.elf" 69632}])
frame_crasher_elf_0002 = frame (4k, fill: [])
frame_goodbye_elf_0000 = frame (4k, fill: [{0 760 CDL_FrameFill_FileData "goodbye.elf" 65536}])
frame_goodbye_elf_0001 = frame (4k, fill: [{0 8 CDL_FrameFill_FileData "goodbye.elf" 69632}])
frame_goodbye_elf_0002 = frame (4k, fill: [])
frame_hello_elf_0000 = frame (4k, fill: [{0 760 CDL_FrameFill_FileData "hello.elf" 65536}])
frame_hello_elf_0001 = frame (4k, fill: [{0 8 CDL_FrameFill_FileData "hello.elf" 69632}])
frame_hello_elf_0002 = frame (4k, fill: [])
frame_monitor_elf_0000 = frame (4k, fill: [{0 4096 CDL_FrameFill_FileData "monitor.elf" 65536}])
frame_monitor_elf_0001 = frame (4k, fill: [{0 3045 CDL_FrameFill_FileData "monitor.elf" 69632}])
frame_monitor_elf_0002 = frame (4k, fill: [{0 8 CDL_FrameFill_FileData "monitor.elf" 73728}])
frame_monitor_elf_0003 = frame (4k, fill: [])
ipcbuf_crasher = frame (4k, fill: [])
ipcbuf_goodbye = frame (4k, fill: [])
ipcbuf_hello = frame (4k, fill: [])
ipcbuf_monitor = frame (4k, fill: [])
monitor_fault_ep = ep
ntfn_crasher = notification
ntfn_goodbye = notification
ntfn_hello = notification
pd_crasher_elf_0001 = pd
pd_goodbye_elf_0001 = pd
pd_hello_elf_0001 = pd
pd_monitor_elf_0001 = pd
pgd_crasher_elf = pgd
pgd_goodbye_elf = pgd
pgd_hello_elf = pgd
pgd_monitor_elf = pgd
pt_crasher_elf_0002 = pt
pt_goodbye_elf_0002 = pt
pt_hello_elf_0002 = pt
pt_monitor_elf_0002 = pt
pud_crasher_elf_0000 = pud
pud_goodbye_elf_0000 = pud
pud_hello_elf_0000 = pud
pud_monitor_elf_0000 = pud
tcb_crasher_elf = tcb (addr: 0x203000,ip: 0x200000,sp: 0x201020,spsr: 0x0,prio: 254,max_prio: 254,affinity: 0,init: [],fault_ep: 0x00000002)
tcb_goodbye_elf = tcb (addr: 0x203000,ip: 0x200000,sp: 0x201020,spsr: 0x0,prio: 254,max_prio: 254,affinity: 0,init: [],fault_ep: 0x00000002)
tcb_hello_elf = tcb (addr: 0x203000,ip: 0x200000,sp: 0x201020,spsr: 0x0,prio: 254,max_prio: 254,affinity: 0,init: [],fault_ep: 0x00000002)
tcb_monitor_elf = tcb (addr: 0x204000,ip: 0x200000,sp: 0x202220,spsr: 0x0,prio: 255,max_prio: 254,affinity: 0,init: [])
}

caps {
cspace_crasher {
0x1: ntfn_crasher (RW)
0x2: monitor_fault_ep (RWGP, badge: 3)
0x3: pgd_crasher_elf
}
cspace_goodbye {
0x1: ntfn_goodbye (RW)
0x2: monitor_fault_ep (RWGP, badge: 2)
0x3: pgd_goodbye_elf
}
cspace_hello {
0x1: ntfn_hello (RW)
0x2: monitor_fault_ep (RWGP, badge: 1)
0x3: pgd_hello_elf
}
cspace_monitor {
0x2: monitor_fault_ep (RW)
0x3: pgd_monitor_elf
}
pd_crasher_elf_0001 {
0x1: pt_crasher_elf_0002
}
pd_goodbye_elf_0001 {
0x1: pt_goodbye_elf_0002
}
pd_hello_elf_0001 {
0x1: pt_hello_elf_0002
}
pd_monitor_elf_0001 {
0x1: pt_monitor_elf_0002
}
pgd_crasher_elf {
0x0: pud_crasher_elf_0000
}
pgd_goodbye_elf {
0x0: pud_goodbye_elf_0000
}
pgd_hello_elf {
0x0: pud_hello_elf_0000
}
pgd_monitor_elf {
0x0: pud_monitor_elf_0000
}
pt_crasher_elf_0002 {
0x0: frame_crasher_elf_0000 (RX)
0x1: frame_crasher_elf_0001 (RW)
0x2: frame_crasher_elf_0002 (RW)
0x3: ipcbuf_crasher (RW)
}
pt_goodbye_elf_0002 {
0x0: frame_goodbye_elf_0000 (RX)
0x1: frame_goodbye_elf_0001 (RW)
0x2: frame_goodbye_elf_0002 (RW)
0x3: ipcbuf_goodbye (RW)
}
pt_hello_elf_0002 {
0x0: frame_hello_elf_0000 (RX)
0x1: frame_hello_elf_0001 (RW)
0x2: frame_hello_elf_0002 (RW)
0x3: ipcbuf_hello (RW)
}
pt_monitor_elf_0002 {
0x0: frame_monitor_elf_0000 (RX)
0x1: frame_monitor_elf_0001 (RX)
0x2: frame_monitor_elf_0002 (RW)
0x3: frame_monitor_elf_0003 (RW)
0x4: ipcbuf_monitor (RW)
}
pud_crasher_elf_0000 {
0x0: pd_crasher_elf_0001
}
pud_goodbye_elf_0000 {
0x0: pd_goodbye_elf_0001
}
pud_hello_elf_0000 {
0x0: pd_hello_elf_0001
}
pud_monitor_elf_0000 {
0x0: pd_monitor_elf_0001
}
tcb_crasher_elf {
cspace: cspace_crasher (guard: 0, guard_size: 56)
fault_ep_slot: monitor_fault_ep (badge: 3,RWGP)
ipc_buffer_slot: ipcbuf_crasher (RW)
vspace: pgd_crasher_elf
}
tcb_goodbye_elf {
cspace: cspace_goodbye (guard: 0, guard_size: 56)
fault_ep_slot: monitor_fault_ep (badge: 2,RWGP)
ipc_buffer_slot: ipcbuf_goodbye (RW)
vspace: pgd_goodbye_elf
}
tcb_hello_elf {
cspace: cspace_hello (guard: 0, guard_size: 56)
fault_ep_slot: monitor_fault_ep (badge: 1,RWGP)
ipc_buffer_slot: ipcbuf_hello (RW)
vspace: pgd_hello_elf
}
tcb_monitor_elf {
cspace: cspace_monitor (guard: 0, guard_size: 56)
ipc_buffer_slot: ipcbuf_monitor (RW)
vspace: pgd_monitor_elf
}
}

irq maps {

}